//*****************************************************************//
//	Testbench for MatrixMultiplication
//	Created By - Vrishbhan Singh Sisodia
//	San Jose State University
//	EE 278
//*****************************************************************//
`timescale 1ns/100ps

module tb;
reg clk_80,rst_80;
reg [8:0] A00_80, A01_80, A02_80, A03_80;
reg [7:0] B00_80, B01_80, B02_80, B03_80;
wire [10:0] AB00_80;

mat_mult m (A00_80, A01_80, A02_80, A03_80, B00_80, B01_80, B02_80, B03_80, 
clk_80, rst_80, AB00_80);

initial begin
	clk_80 = 1'b0;
	repeat (1000) clk_80 = #5 ~clk_80;
	//$finish;
end
initial begin
		rst_80 = 1'b1;
		#10
		rst_80 = 1'b0;
end

initial begin
	A00_80 = 0;
	B00_80 =  0;
	A01_80 = 0;
	B01_80 = 0;
	A02_80 = 0;
	B02_80 = 0;
	A03_80 = 0;
	B03_80 = 0;
	#5;
	A00_80 = 10;//X00
	A01_80 = 20;//X01
	A02_80 = 30;//X02
	A03_80 = 40;//X03
	#0;
	B00_80 =  13;//Y00 = 0.1
	B01_80 = 77;//Y10 = 0.6
	B02_80 = 102;//Y20 = 0.8
	B03_80 = 205;//Y20 = -0.4
	#10;
	B00_80 =  26;//Y01 = 0.2
	B01_80 = 166;//Y11 = -0.7
	B02_80 = 90;//Y21 = 0.7
	B03_80 = 38;//Y31 = 0.3
	#10;
	B00_80 =  38;//Y02 = 0.3
	B01_80 = 154;//Y12 = -0.8
	B02_80 = 77;//Y22 = 0.6
	B03_80 = 230;//Y32 = -0.2
	#10;
	B00_80 =  192;//Y03 = -0.5
	B01_80 = 115;//Y13 = 0.9
	B02_80 = 64;//Y23 = 0.5
	B03_80 = 13;//Y33 = 0.1
	#10;
	A00_80 = 50;//X10
	A01_80 = 60;//X11
	A02_80 = 70;//X12
	A03_80 = 80;//X13
	#0;
	B00_80 =  13;//Y00 = 0.1
	B01_80 = 77;//Y10 = 0.6
	B02_80 = 102;//Y20 = 0.8
	B03_80 = 205;//Y20 = -0.4
	#10;
	B00_80 =  26;//Y01 = 0.2
	B01_80 = 166;//Y11 = -0.7
	B02_80 = 90;//Y21 = 0.7
	B03_80 = 38;//Y31 = 0.3
	#10;
	B00_80 =  38;//Y02 = 0.3
	B01_80 = 154;//Y12 = -0.8
	B02_80 = 77;//Y22 = 0.6
	B03_80 = 230;//Y32 = -0.2
	#10;
	B00_80 =  192;//Y03 = -0.5
	B01_80 = 115;//Y13 = 0.9
	B02_80 = 64;//Y23 = 0.5
	B03_80 = 13;//Y33 = 0.1
	#10;
	A00_80 = 90;//X20
	A01_80 = 100;//X21
	A02_80 = 110;//X22
	A03_80 = 120;//X23
	#0;
	B00_80 =  13;//Y00 = 0.1
	B01_80 = 77;//Y10 = 0.6
	B02_80 = 102;//Y20 = 0.8
	B03_80 = 205;//Y20 = -0.4
	#10;
	B00_80 =  26;//Y01 = 0.2
	B01_80 = 166;//Y11 = -0.7
	B02_80 = 90;//Y21 = 0.7
	B03_80 = 38;//Y31 = 0.3
	#10;
	B00_80 =  38;//Y02 = 0.3
	B01_80 = 154;//Y12 = -0.8
	B02_80 = 77;//Y22 = 0.6
	B03_80 = 230;//Y32 = -0.2
	#10;
	B00_80 =  192;//Y03 = -0.5
	B01_80 = 115;//Y13 = 0.9
	B02_80 = 64;//Y23 = 0.5
	B03_80 = 13;//Y33 = 0.1
	#10;
	A00_80 = 130;//X30
	A01_80 = 140;//X31
	A02_80 = 150;//X32
	A03_80 = 160;//X33
	#0;
	B00_80 =  13;//Y00 = 0.1
	B01_80 = 77;//Y10 = 0.6
	B02_80 = 102;//Y20 = 0.8
	B03_80 = 205;//Y20 = -0.4
	#10;
	B00_80 =  26;//Y01 = 0.2
	B01_80 = 166;//Y11 = -0.7
	B02_80 = 90;//Y21 = 0.7
	B03_80 = 38;//Y31 = 0.3
	#10;
	B00_80 =  38;//Y02 = 0.3
	B01_80 = 154;//Y12 = -0.8
	B02_80 = 77;//Y22 = 0.6
	B03_80 = 230;//Y32 = -0.2
	#10;
	B00_80 =  192;//Y03 = -0.5
	B01_80 = 115;//Y13 = 0.9
	B02_80 = 64;//Y23 = 0.5
	B03_80 = 13;//Y33 = 0.1
	#20;
	$finish;
end

endmodule